// stage1
module stage1
	(
		assign 
	);
)
