// stage1
module stage1
	(
		assign always_comb begin
			
		end
	);

endmodule
