// stage1
module stage1(CLOCK_50, SW, KEY);
	input CLOCK_50;
	input [9:0] SW;
	input [3:0] KEY;

	contorl c0();

	datapath d0();



endmodule

module control();

endmodule

module datapath();

endmodule
//  RAM 64 words x 32 bits
