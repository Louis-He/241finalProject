// stage1
module stage1(CLOCK_50, SW, KEY);
	input CLOCK_50;
	input [9:0] SW;
	input [3:0] KEY;
endmodule

module control();

endmodule

module datapath();

endmodule
